//
//
//---- Top entity
module top (
 input  ICE_PB,
 output LED_R
);
 wire w0;
 assign ICE_PB = w0;
 assign w0 = LED_R;
endmodule

